`timescale 1ns / 1ps


module Adder_Nbit(
    input [31:0] A,
    input [31:0] B,
    output [31:0] C
    );
    assign C = A + B;
endmodule
